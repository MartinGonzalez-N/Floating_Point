`define PIPLINE